//////////////////////////////////////////MUX_2_1_MODULE/////////////////////////////////////////////////////
module mux2_1(input [31:0] ina,inb, input sel, 
              output [31:0] out);

endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////PC_MODULE///////////////////////////////////////////////////////////////
module PC(input clk,res,write, 
          input [31:0] in, 
          output reg [31:0] out);
  
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////INSTRUCTION_MEMORY/////////////////////////////////////////////////////
module instruction_memory(input [9:0] address, 
                          output reg[31:0] instruction);

  reg [31:0] codeMemory [0:1023];
  
  initial $readmemh("code.mem", codeMemory);

endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////ADDER_MODULE//////////////////////////////////////////////////////
module adder(input [31:0] ina,inb, 
             output reg[31:0] out);

endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////



//////////////////////////////////////////////IF//////////////////////////////////////////////////////////////
module IF (input clk,reset,PCSrc,PC_write, 
           input [31:0] PC_Branch, 
           output [31:0] PC_IF, INSTRUCTION_IF)

endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////



///////////////////////////////////REGISTER_FILE_MODULE///////////////////////////////////////////////////////
module registers(input clk,reg_write,
                 input [4:0] read_reg1,read_reg2,write_reg,
                 input [31:0] write_data,
                 output [31:0] read_data1,read_data2);

endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////



//////////////////////////////////////////IMM_GEN_MODULE/////////////////////////////////////////////////////
module imm_gen(input [31:0] in,
               output reg [31:0] out);
  
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////



//////////////////////////////////////////////ID_MODULE////////////////////////////////////////////////////////
module ID(input clk,
          input [31:0] PC_ID,INSTRUCTION_ID,
          input RegWrite_WB,
          input [31:0] ALU_DATA_WB,
          input [4:0] RD_WB,
          output [31:0] IMM_ID,
          output [31:0] REG_DATA1_ID,REG_DATA2_ID,
          output [2:0] FUNCT3_ID,
          output [6:0] FUNCT7_ID.
          output [6:0] OPCODE_ID
          output [4:0] RD_ID,
          output [4:0] RS1_ID,
          output [4:0] RS2_ID);
  
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////



////////////////////////////////////////PIPELINE_REG_MODULES///////////////////////////////////////////////////
module IF_ID_reg(input clk,reset,write,
                 input [31:0] pc_in,instruction_in
                 ouput reg [31:0] pc_out,instruction_out);
  
endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////



/////////////////////////////////////////////RISC_V_IF_ID/////////////////////////////////////////////////////
module RISC_V_IF_ID(input clk,reset,
                    input IF_ID_write, PCSrc, PC_write,
                    input [31:0] PC_Branch,
                    input RegWrite_WB,
                    input [31:0] ALU_DATA_WB,
                    input [4:0] RD_WB,
                    output [31:0] PC_ID, INSTRUCTION_ID, IMM_ID, REG_DATA1_ID, REG_DATA2_ID
                    output [2:0] FUNCT3_ID,
                    output [6:0] FUNCT7_ID, OPCODE_ID,
                    output [4:0] RD_ID, RS1_ID, RS2_ID);


endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////
